package msnw_pkg;

// Import the UVM class library  and UVM automation macros
 import uvm_pkg::*;
`include "uvm_macros.svh"
`include "msnw_trans.sv"
`include "msnw_err_trans.sv"
`include "msnw_monitor.sv"
`include "msnw_in_driver.sv"
`include "msnw_out_driver.sv"
`include "msnw_sequencer.sv"
`include "msnw_agent.sv"
//  `include "msnw_scoreboard.sv"
`include "msnw_env.sv"

endpackage : msnw_pkg

